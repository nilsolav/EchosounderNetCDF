netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
    :title = "Echogram scrutiny masks";
	
group: Interpretation {
	group: v1 { // subsequent versions of this interpretation get put in new subgroups, using the numbering system v1, v2, etc.
		// SUGGESTIONS OF THINGS TO ADD:
		// - consider a separate implementation of layers, as per LSSS
		// - link to categorisation database and database version
		// - name of echosounder files that the data came from??
		
		:version = "1"; // increasing integers
		:version_save_date = "20190903T154023Z"; // ISO8601 format
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		
		types:
			// Note: empty_water == LSSS erased; no_data == LSSS excluded
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			// Storing 3D regions is not yet done, but we include the region dimension here anyway
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t; // ragged array for region ping times
		dimensions:
			regions = 3; // varies to suit data. Could also be unlimited
			channels = 3; // varies to suit data
			categories = 5; // varies to suit data.
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
				
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			// simple example regions
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  0.0, 20.5, 55.0;
			max_depth = 10.0, 42.0, 125.2;
			start_time = 13189164120001, 13189164121000, 13189164124000;
			end_time =   13189164123004, 13189164124000, 13189164131000;
			region_id = 1, 5, 234;
			region_name = "region1", "region2", "";
			region_provenance = "KORONA-2.6.0;LSSS", "Echoview - template ABC", "Manual inspection";
			region_comment = "", "", "whale!";
			region_category_names = "herring", "krill", "seal", "lion", "platypus";
			region_category_proportions = 0.9, 0.1, 0.45, 0.40, 0.10;
			region_category_ids = 1, 1, 234, 234, 234;
			region_type = analysis, empty_water, analysis;
			channel_names = "18kHz WBT ABC", "38kHz WBT ZYX", "120kHz GPT 123";
			region_channels = 5, 7, 7;
			mask_times = {13189164120001, 13189164121002, 13189164122003, 13189164123004}, 
						 {13189164121000, 13189164122000, 13189164123000, 13189164124000}, 
						 {13189164124000, 13189164125000, 13189164126000, 13189164127000, 13189164128000, 13189164129000, 13189164131000};
			mask_depths = {{0.0, 5.0}, {0.0, 4.0, 5.0, 10.0}, {0.0, 10.0}, {0.0, 10.0}}, {{20.5, 25.0}, {30.5, 35.0}, {35.5, 40.0}, {40.0, 42.0}}, {{55.0, 105.0}, {60.0, 80.2, 100.6, 115.0}, {55.0, 107.0}, {55.0, 110.0}, {55.0, 115.6}, {55.0, 125.2}, {60, 115}};
		}
	}
}
