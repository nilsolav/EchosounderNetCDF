netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
    :title = "Echogram scrutiny masks";
	
group: Interpretation {
	// SUGGESTIONS OF THINGS TO ADD:
	// - consider a separate implementation of layers, as per LSSS
	// - link to categorisation database and database version
	// - name of echosounder files that the data came from??
	
	types:
		// Note: empty_water == LSSS erased; no_data == LSSS excluded
		byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
		// Storing 3D regions is not yet done, but we include the region dimension here anyway
		byte enum region_dim_t {twoD = 0, threeD = 1};
		float(*) mask_depth_t;
		uint64(*) mask_time_t;
	dimensions:
		regions = 3; // varies to suit data. Could also be unlimited
		channels = 3; // varies to suit data
	variables:
		float sound_speed;
			sound_speed:long_name = "Sound speed used to convert echo time into range";
			sound_speed:standard_name = "speed_of_sound_in_sea_water";
			sound_speed:units = "m/s";
			sound_speed:valid_min = 0.0;

		// The bounding box of each region
		float min_depth(regions);
			min_depth:long_name = "Minimum depth for each region";
			min_depth:units = "m";
			min_depth:valid_min = 0.0;
		float max_depth(regions);
			max_depth:long_name = "Maximum depth for each regions";
			max_depth:units = "m";
			max_depth:valid_min = 0.0;
		uint64 start_time(regions);
			start_time:long_name = "Timestamp of the earliest data point in each region";
			start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
			start_time:axis = "T";
			start_time:calendar = "gregorian";
			start_time:standard_name = "time";
		uint64 end_time(regions);
			end_time:long_name = "Timestamp of the latest data point in each region";
			end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
			end_time:axis = "T";
			end_time:calendar = "gregorian";
			end_time:standard_name = "time";
			
		region_dim_t region_dimension; 
			region_dimension:long_name = "Region dimension";

		int id(regions);
			id:long_name = "Dataset-unique identification number for each region";
		string name(regions);
			name:long_name = "Name of each region";
		string provenance(regions);
			provenance:long_name = "Provenance of each region"; 
		string comment(regions);
			comment:long_name = "Comment for each region";
		string category(regions);
			category:long_name = "Categorisation for each region";
		region_t region_type(regions);
			region_type:long_name = "Region type";
		
		string channel_names(channels);
			channel_names:long_name = "Echosounder channel names";
		uint region_channels(regions);
			region_channels:long_name = "Echosounder channels that this region applies to";
			region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
			region_channels:_FillValue = 4294967295; // 2^32-1
			
		mask_time_t mask_times(regions);
			mask_times:long_name = "Timestamp of each mask point";
			mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
			mask_times:axis = "T";
			mask_times:calendar = "gregorian";
			mask_times:standard_name = "time";
		mask_depth_t mask_depths(regions);
			mask_depths:long_name = "Depth pairs of mask";
			mask_depths:units = "m";
			mask_depths:valid_min = 0.0;
	
	data:
	    // simple example regions
		region_dimension = twoD;
		sound_speed = 1496;
		min_depth =  0.0, 20.5, 55.0;
		max_depth = 10.0, 42.0, 125.2;
		start_time = 13210680841000, 13210680843000, 13210680845000;
		end_time =   13210680847000, 13210680846000, 13210680850000;
		id = 1, 5, 234;
		name = "region1", "region2", "";
		provenance = "KORONA-2.6.0;LSSS", "Echoview - template ABC", "Manual inspection";
		comment = "", "", "whale!";
		category = "herring", "", "whale";
		region_type = analysis, empty_water, analysis;
		channel_names = "18kHz WBT ABC", "38kHz WBT ZYX", "120kHz GPT 123";
		region_channels = 5, 7, 7;
		mask_times = {13210680841000, 13210680842000, 13210680843000, 13210680847000}, 
		             {13210680843000, 13210680844000, 13210680845000, 13210680846000}, 
					 {13210680845000, 13210680846000, 13210680846000, 13210680847000, 13210680848000, 13210680849000, 13210680850000};
		mask_depths = {0.0, 5.0, 0.0, 8.0, 0.0, 10.0, 0.0, 10.0}, {20.5, 25.0, 30.5, 35.0, 35.5, 40.0, 40.0, 42.0}, {55.0, 105.0, 60.0, 80.2, 100.6, 115.0, 55.0, 107.0, 55.0, 110.0, 55.0, 115.6, 55.0, 125.2};	
	}
}
